library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity pacman_game is
   Port (
		clk       : in  STD_LOGIC
--      reset     : in  STD_LOGIC;
--      vga_HS    : out STD_LOGIC;
--      vga_VS    : out STD_LOGIC;
--      pixel_x   : out INTEGER range 0 to 1279;
--      pixel_y   : out INTEGER range 0 to 1023
--		  
--      --PIXEL_COLOR : out STD_LOGIC_VECTOR(11 downto 0)
   );
end pacman_game;

architecture Behavioral of pacman_game is



begin
	
end Behavioral;