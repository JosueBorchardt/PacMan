library verilog;
use verilog.vl_types.all;
entity video_controller_vlg_vec_tst is
end video_controller_vlg_vec_tst;
